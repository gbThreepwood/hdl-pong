`default_nettype none



module vga_test_pattern_generator #(
    parameter c_COLOR_BIT_WIDTH = 3,
    parameter c_VISIBLE_COLUMNS = 640,
    parameter c_VISIBLE_ROWS = 480,
    parameter c_TOTAL_COLUMNS = 800,
    parameter c_TOTAL_ROWS = 525
)
(
    input wire i_Clk,
    input wire [3:0] i_PatternSelect,
    input wire i_HSync,
    input wire i_VSync,
    input wire [9:0] i_ColCount,
    input wire [9:0] i_RowCount,
    output wire o_HSync,
    output wire o_VSync,
    output reg [c_COLOR_BIT_WIDTH - 1:0] o_VideoRed = 0,
    output reg [c_COLOR_BIT_WIDTH - 1:0] o_VideoGreen = 0,
    output reg [c_COLOR_BIT_WIDTH - 1:0] o_VideoBlue = 0
);

    assign o_HSync = i_HSync;
    assign o_VSync = i_VSync;

    // Declare 3 bit wide (by default) arrays with a depth of 16 for each of the three colors
    // I.e. we have sixteen three bit wide arrays for each color
    // The patterns are generated by changing the 3-bit value depending on the current row and
    // column counter value.
    wire [c_COLOR_BIT_WIDTH - 1:0] RedPattern [0:15];
    wire [c_COLOR_BIT_WIDTH - 1:0] GreenPattern [0:15];
    wire [c_COLOR_BIT_WIDTH - 1:0] BluePattern [0:15];

    assign RedPattern   [0] = 0;
    assign GreenPattern [0] = 0;
    assign BluePattern  [0] = 0;

    assign RedPattern   [1] = (i_ColCount < c_VISIBLE_COLUMNS && i_RowCount < c_VISIBLE_ROWS) ? { c_COLOR_BIT_WIDTH{1'b1} } : 0;
    assign GreenPattern [1] = 0;
    assign BluePattern  [1] = 0;

    assign RedPattern   [2] = 0;
    assign GreenPattern [2] = (i_ColCount < c_VISIBLE_COLUMNS && i_RowCount < c_VISIBLE_ROWS) ? { c_COLOR_BIT_WIDTH{1'b1} } : 0;
    assign BluePattern  [2] = 0;

    assign RedPattern   [3] = 0;
    assign GreenPattern [3] = 0;
    assign BluePattern  [3] = (i_ColCount < c_VISIBLE_COLUMNS && i_RowCount < c_VISIBLE_ROWS) ? { c_COLOR_BIT_WIDTH{1'b1} } : 0;

    // Chessboard pattern
    assign RedPattern   [4] = i_ColCount[5] ^ i_RowCount[5] ? {c_COLOR_BIT_WIDTH{1'b1}} : 0;
    assign GreenPattern [4] = RedPattern[4];
    assign BluePattern  [4] = RedPattern[4];


    // Split the display in to 8 color bars

    wire [6:0] w_BarWidth;
    wire [3:0] w_BarSelect;

    assign w_BarWidth = c_VISIBLE_COLUMNS / 8;

    assign w_BarSelect = i_ColCount < w_BarWidth*1 ? 0 :
                         i_ColCount < w_BarWidth*2 ? 1 :
                         i_ColCount < w_BarWidth*3 ? 2 :
                         i_ColCount < w_BarWidth*4 ? 3 :
                         i_ColCount < w_BarWidth*5 ? 4 :
                         i_ColCount < w_BarWidth*6 ? 5 :
                         i_ColCount < w_BarWidth*7 ? 6 :
                         i_ColCount < w_BarWidth*8 ? 7 : 8;
    
    assign RedPattern   [5] = w_BarSelect[2] ? {c_COLOR_BIT_WIDTH{1'b1}} : 0; //w_BarSelect > 3 ? 1 : 0;
    assign GreenPattern [5] = w_BarSelect[1] ? {c_COLOR_BIT_WIDTH{1'b1}} : 0;
    assign BluePattern  [5] = w_BarSelect[0] ? {c_COLOR_BIT_WIDTH{1'b1}} : 0;

    // Generate some colors
    reg [2:0] r_RedPattern = 0;
    reg [2:0] r_GreenPattern = 0;
    reg [2:0] r_BluePattern = 0;

    assign RedPattern   [6] = r_RedPattern;
    assign GreenPattern [6] = r_GreenPattern;
    assign BluePattern  [6] = r_BluePattern;

    always @(posedge i_Clk) begin
 
        if (i_ColCount < c_VISIBLE_COLUMNS && i_RowCount < c_VISIBLE_ROWS) begin
            
            if (i_ColCount <= 160) begin
                r_RedPattern    <= 3'b111;
                r_GreenPattern  <= 3'b000;
                r_BluePattern   <= 3'b000;
            end
            else if ((i_ColCount > 160) && (i_ColCount < 320)) begin
                r_RedPattern    <= 3'b000;
                r_GreenPattern  <= 3'b111;
                r_BluePattern   <= 3'b000;
            end
            else begin
                r_RedPattern    <= 3'b000;
                r_GreenPattern  <= 3'b000;
                r_BluePattern   <= 3'b111;
            end
        end
        else begin
            r_RedPattern    <= 3'b000;
            r_GreenPattern  <= 3'b000;
            r_BluePattern   <= 3'b000;           
        end
    end


    // Read a bitmap
    reg [12:0] r_pixel_addr = 0;
    wire [8:0] w_pixel_data;

    always @(posedge i_Clk) begin

        if (i_ColCount < c_VISIBLE_COLUMNS && i_RowCount < c_VISIBLE_ROWS) begin
            r_pixel_addr <= i_ColCount + (i_RowCount * 160);
        end
        else begin
            r_pixel_addr <= 0;
        end

    end

    block_ram #(
        .ADDR_WIDTH(13), // We need to address 4800 9-bit values
        .DATA_WIDTH(9),  // Each memory location should hold 3x3 bit of color information
        .MEM_INIT_FILE("test_image.mem")
    ) bitmap_block_ram_inst
    (
        .i_clk(i_Clk),
        .i_write_en(1'b0),
        .i_addr(r_pixel_addr),
        .i_din(),
        .o_dout(w_pixel_data)
    );

    // Read a bitmap from block RAM
    assign RedPattern   [7] = w_pixel_data[2:0];
    assign GreenPattern [7] = w_pixel_data[5:3];
    assign BluePattern  [7] = w_pixel_data[8:6];


    // Line drawing algorithm test
    assign RedPattern   [0] = 0;
    assign GreenPattern [0] = 0;
    assign BluePattern  [0] = 0;


    always @(posedge i_Clk) begin
        case (i_PatternSelect)
            4'h0: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
            4'h1: begin
                o_VideoRed   <= RedPattern   [1];
                o_VideoGreen <= GreenPattern [1];
                o_VideoBlue  <= BluePattern  [1];
            end
            4'h2: begin
                o_VideoRed   <= RedPattern   [2];
                o_VideoGreen <= GreenPattern [2];
                o_VideoBlue  <= BluePattern  [2];
            end
            4'h3: begin
                o_VideoRed   <= RedPattern   [3];
                o_VideoGreen <= GreenPattern [3];
                o_VideoBlue  <= BluePattern  [3];
            end
            4'h4: begin
                o_VideoRed   <= RedPattern   [4];
                o_VideoGreen <= GreenPattern [4];
                o_VideoBlue  <= BluePattern  [4];
            end
            4'h5: begin
                o_VideoRed   <= RedPattern   [5];
                o_VideoGreen <= GreenPattern [5];
                o_VideoBlue  <= BluePattern  [5];
            end
            4'h6: begin
                o_VideoRed   <= RedPattern   [6];
                o_VideoGreen <= GreenPattern [6];
                o_VideoBlue  <= BluePattern  [6];
            end
            4'h7: begin
                o_VideoRed   <= RedPattern   [7];
                o_VideoGreen <= GreenPattern [7];
                o_VideoBlue  <= BluePattern  [7];
            end
            4'h8: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
            4'h9: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
            4'hA: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
            4'hB: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
            4'hC: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
            4'hD: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
            4'hE: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
            4'hF: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
            default: begin
                o_VideoRed   <= RedPattern   [0];
                o_VideoGreen <= GreenPattern [0];
                o_VideoBlue  <= BluePattern  [0];
            end
        endcase
    end

endmodule
