`default_nettype none

module encoder_read();

endmodule
